`include "alu.sv"

module top (
  input  logic clk,
  output logic out
);

alu DUT();

endmodule