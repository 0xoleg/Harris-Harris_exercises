`include "exercise5.12/tb5.12.sv"

module top (
  input  logic clk,
  output logic out
);

//testbench tb();

endmodule